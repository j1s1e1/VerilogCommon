module Precision();
// This file just hides all the other files in these folders
// Since some FPGA software does not use folders in design sources

add();
abs();
add_matrix();
delay_v();
divide_vector();
divide_vector_by_scalar();
exponent();
min_index_matrix_row();
min_vector();
multiply_vector();
set_value();
subtract();
subtract_scalar_from_vector();
subtract_vector();
sum_vector();
two_int_power();

half_max_v();
half_min_v();
half_max_abs_v();
half_integer_part();

fixed_add();
fixed_divide();
fixed_multiply();
fixed_integer_part();
fixed_two_int_power();

single_integer_part();
single_max_abs();
single_max_v();

endmodule