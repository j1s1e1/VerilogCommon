`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/02/2020 04:59:41 PM
// Design Name: 
// Module Name: half_base2_exp
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module half_base2_exp
(
input clk,
input in_valid,
input [15:0] a,
output logic out_valid,
output logic [15:0] c
);



endmodule
